module UART_Control(
		input           Clk             , // Clock
		input           Rst_n           , // Reset
		input	[47:0]	 x_coord         ,
		input [47:0]    y_coord         ,
		input [47:0]    z_coord         ,
		output          Tx                // RS232 TX line.
	);
	
/////////////////////////////////////////////////////////////////////////////////////////
reg [7:0]    	TxData     	; // Data to transmit.
wire          	TxDone          ; // Trnasmission completed. Data sent.
wire            tick		; // Baud rate clock
reg          	TxEn            ;
wire [3:0]      NBits    	;
wire [15:0]    	BaudRate        ; //328; 162 etc... (Read comment in baud rate generator file)

/////////////////////////////////////////////////////////////////////////////////////////
assign 		BaudRate = 16'd325; 	//baud rate set to 9600 for the HC-06 bluetooth module. Why 325? (Read comment in baud rate generator file)
assign 		NBits = 4'b1000	;	//We send/receive 8 bits
/////////////////////////////////////////////////////////////////////////////////////////


//Make connections between Tx module and TOP inputs and outputs and the other modules
UART_rs232_tx I_RS232TX(
   	.Clk(Clk)            	,
    	.Rst_n(Rst_n)         	,
    	.TxEn(TxEn)           	,
    	.TxData(TxData)      	,
   	.TxDone(TxDone)      	,
   	.Tx(Tx)               	,
   	.Tick(tick)           	,
   	.NBits(NBits)
    );

//Make connections between tick generator module and TOP inputs and outputs and the other modules
UART_BaudRate_generator I_BAUDGEN(
    	.Clk(Clk)               ,
    	.Rst_n(Rst_n)           ,
    	.Tick(tick)             ,
    	.BaudRate(BaudRate)
    );


wire [7:0]str[0:61];

assign str[0]=8'h44;//D
assign str[1]=8'h65;//E
assign str[2]=8'h73;//S
assign str[3]=8'h69;//I
assign str[4]=8'h72;//R
assign str[5]=8'h65;//E
assign str[6]=8'h64;//D
assign str[7]=8'h20;
assign str[8]=8'h73;//S
assign str[9]=8'h6F;//O
assign str[10]=8'h75;//U
assign str[11]=8'h6E;//N
assign str[12]=8'h64;//D
assign str[13]=8'h20;
assign str[14]=8'h64;//D
assign str[15]=8'h65;//E
assign str[16]=8'h74;//T
assign str[17]=8'h65;//E
assign str[18]=8'h63;//C
assign str[19]=8'h74;//T
assign str[20]=8'h65;//E
assign str[21]=8'h64;//D
assign str[22]=8'h21;//!
assign str[23]=8'h21;//!
assign str[24]=8'h20;
assign str[25]=8'h0A;
assign str[26]=8'h43;//C
assign str[27]=8'h6F;//O
assign str[28]=8'h6F;//O
assign str[29]=8'h72;//R
assign str[30]=8'h64;//D
assign str[31]=8'h73;//S
assign str[32]=8'h3A;//:
assign str[33]=8'h0A;
assign str[34]=8'h58;//X
assign str[35]=8'h3A;//:

assign str[36]=x_coord[47:40];//
assign str[37]=x_coord[39:32];//
assign str[38]=x_coord[31:24];//
assign str[39]=x_coord[23:16];//
assign str[40]=x_coord[15:8];//
assign str[41]=x_coord[7:0];//

assign str[42]=8'h0A;
assign str[43]=8'h59;//Y
assign str[44]=8'h3A;//:

assign str[45]=y_coord[47:40];//
assign str[46]=y_coord[39:32];//
assign str[47]=y_coord[31:24];//:
assign str[48]=y_coord[23:16];//:
assign str[49]=y_coord[15:8];//:
assign str[50]=y_coord[7:0];//:

assign str[51]=8'h0A;
assign str[52]=8'h5A;//Z
assign str[53]=8'h3A;//:

assign str[54]=z_coord[47:40];//
assign str[55]=z_coord[39:32];//
assign str[56]=z_coord[31:24];//
assign str[57]=z_coord[23:16];//
assign str[58]=z_coord[15:8];//
assign str[59]=z_coord[7:0];//

assign str[60]=8'h0A;
assign str[61]=8'h0A;

parameter s0=0,s1=1,s2=2,s3=3;
reg [1:0]current_state;
reg [1:0]next_state;
reg [5:0] n=0;
integer N=61;


always@(posedge tick or negedge Rst_n) begin
	if (~Rst_n) begin
		current_state <= s3;
	end
	else
		current_state <= next_state;
end

always@(posedge tick)begin
	case(current_state)
		s0: begin		
			TxEn<=0;
			TxData <= str[n];
			next_state <= s1;
		end
		s1: begin
			TxEn<=1;
			next_state <= s2;
		end
		s2: begin
			if(TxDone) begin
				TxEn <= 0;
				if (n<N) begin
					n = n + 1;
					next_state<=s0;
				end
			end
		end
		s3: begin
			n=0;
			next_state <= s0;
		end
	endcase
end


endmodule
